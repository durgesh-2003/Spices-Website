���� JFIF       �� .Exif  MM *    @      M  @            �� C 
	
		
$ &%# #"(-90(*6+"#2D26;=@@@&0FKE>J9?@=�� C=)#)==================================================�� 
�" ��           	
�� �   } !1AQa"q2���#B��R��$3br�	
%&'()*456789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz���������������������������������������������������������������������������        	
�� �  w !1AQaq"2�B����	#3R�br�
$4�%�&'()*56789:CDEFGHIJSTUVWXYZcdefghijstuvwxyz��������������������������������������������������������������������������   ? 񞦵,�%�⳸�m�A���=���veV�"�yj���{W[ix��jW�;��eIj|�ƦN��\�F�g���7l��)@frI��*	Š�.�G��Qʢ��'�pj�����v� n��[��*HF���R?�hO&���x<�in$�%���	�㧽es{[B�ď�^�}���Z4��V>Yde����������mVx�w�R�\�H��}�q�VD�r�z����<��.b@˒r{�lt�뚬qk�vki.lci@��#����f������0��SV�ԯ�-��1ǐn�k��4�,YhRjqMke<Y�%�]������Su-J='U���4�+c��g�Fp0F	<��:��ki�4q[i"y���2H�לS颷p�v��h��]�zz�\X��d�d�dl}ާ ��d�Uo���#\}`Ɨ�"8� 0x�<q���l_x�t��D�Y��,A1��l;c�$��\Ϳ�/5Rɵ)���$33o�О��O�	+�Bm��[}0͡�N��YKj��i��@��qV�ۻ����O����{E�P>|�}���E7W���<W#��Q��Y|�pdW z�*ĚL7��i� �P�����]B�+�����hz��i�+Km�j�v�w7�gm1���e�zu9>�GJ��4k�Z-׮�8$S�U�p`x���i��[�x�b��(��˿�w�3�diZuĂmB�/2+&1t��<g뎔լŪjۖ�|GuqkcdaC�&�m<���8��}fk��=�Y�OG�R#��=x�ָ�W��.5Z�0ƍ�%�q�Υ�n,�t+;�s4ڻ92�n��a��RI�Td��z���#(Om��y�ͨ��]2 Bά��κ�jm���L�/�k����U�u`Lv�Ќ�m��/#}�G/5�'g�W�R���!@8�f�����b�Rۑ�� <�k��t��4�K=ζ=G1ݐ� �� ^�a�2;��.種F+�XA��p�� ?�jY]��1+��[ӑ���U��^�\*ju"F����HF�<t�Ӑ'�Nd	�i�=?3T�x��"��>���V�-�'b���	���^kVv�o�3|ݓ�-%�a\�-�1�|��U'̺ͬQe� ���?�	�b�E�N���_�n<0V���y�u��.%�y$�B�ʫ ~i������褝�����jKr�+�8��tf8�?�eI<�]��6C+5���|���Qr�_�R۩V�[	�V8����J�p#��k�ك�++�V9�>�~<WE*v�{؉I�ū4��V�f_7-��H�rq�zO��D���{Fah\�F��s��5���Ĉ�E� ,� 2�S�º��'���7���͐� .?����q�֟3�n�۝׏tv�|1l���?60;�s���Ƽ7�W�g�;WL0��#<0�}+p�P�ϭ|�i�E��-��;�S���~�Wrz4p�Z&'��d�f�BLR�q����U����{q���h@?S[�6R�n�#(�������s�w-�k�qLv�de��� �҃N3����|�����>4��	�O^j�ɚK+-P �� >��oʹ�Ks�#kcf ��ۦ��]E���<�q%�.�X�=>��>V����M���[ٍ*;�$u0|�=29�s:��^�_����C{��6��0Ǡ��W=#�B��-Fr;�qI�G%�U��6il��'��
ґ��±�ڴ���%0�����mﶈ6�l�dtz���P�w��K�OܡbO}�����Y��gR�����I���&W������5��&��������x#?��]����G�2��UNP}}8�}�'��5h�Bg�A�N	Ϯ=8��Д�^���Iom{g&S�Ł���qUݴ�f)f��H��	Ϧ*ƛp"���=6��'S�A�SW�9z4Oy��2J�V%a��C�|d~4��nۊ�X/�n-J-��I�y2H7}{��nLפH�2��y鏭Y�/���6ב� �y���A}$���ZD1�ªG֜tKMX��}� ��r+������E���2� �\���Բ�Fp{��ѵ���7O���:��D�*�Sz����:��I�|�rOp�v<��jiW-y��<�4E��#����(��X�$�W?�Դ8O���^����?�roQ�}B�k�:�g������b ��
銲��9sJ��d�� �#P=���TL�Q�
�[yf����YSko����Ti���\"�X��f���ZII� 0&�I�8�kI��A����G�KC��N~��2H9��Q�x���p�TrXJ3�kc����L��% ���5v���|�J�U�k[���?:�t�ّ�@�WK Α�b��C�ں襸�[���K�saP�מk����;�p��R�y��hSOi1��(n��3t� ��N8%���Q=ʦ]Ӵ�5;���C���rYW�ϱ�t��~�{�;�.,b��	%a����=�N
��9���w��ۇ��`ܹ��^�p)��x������:42J�<F��$�ӜT[]Mo}�.���̰D����4�*N�s��%�u����ZCd��K{1��S�Ǳ?�-��z�JK�����$�R�6O�����+k�'N���t>Kۇ��$�~b��8=�Il�iu,����zdBA�<����ٻ���X��hj��o��)4��
[��V�G<V����ؠ��%���Y#�� �\�9q��=��oai����"��.m�/)b z���J���ˑ�$^(�tk��t�	"�L0P���r?��Z_��]h�^����d \��=zv��cM�����o삙e�,���I<��Yri�Z�ޫ��%����.OLz��U�웻�mɏX��\�]�"b��lI�>)���xB�d�����U}��R�Qh������DX�8HR��_PO㊣s�Y�Yi��^+-��$�s�s��N���4|-z�=֣u�mmq�/0�\��I���}�mB�3k�"q�ʏ��9��jֽym>�2�㱃�NN�׽Aix�F�m�����:p�F�M]Z����<�xi/l-��x���a����A��UkP��K�K8lg*�f�n珓�d��VU�I��]M�k���Di�V�YGN�[ն�˒ʛ�`e�}9���]��%s��͢� h�;����<��k��4{��h�`�^sd���/����x�a`�_v����ֽ3&k[�csr{VR����nǋji�]�ш����j�JU�V
}Oj��EehI�ᑀ�9��P�����Zjg�^����X�zWA��CY�v$31;������	rz��_��h%V�8=c^�4ZEҫ���*β M���������p�F��Ϯs�W#�].7J����3��E���#�EU�A��u�:��֢�#ӧ+�i-~߲�7�Q�<r��~5��q4�$�,J�p �lr>��ާ��k�6��!T;Fv���g�r�_�o�'KxDP�Vd6�ݎ:8�E*4�[��h95y�m���P�O-~��F��N=	8:
Ľ�I6�����T�.�y����sZ� ��i��~���!U�ݟ�����\��ҙ���F�,#�ݿ 9�޽J���9j6���F�{7T
��FJ��˃�V��t"���̋'�!���˧��9$s�ZC#FJ������������ 2�� N8�����E%t��l��%���H�w#�C\��/y�x��Z�X�c�Q�k����W�5�V�]C����򿉯u�����.�g߸		��k�۹�R3i�}�K-Ab��M�E�!$S���?㌉���$��ۨ� �w���a��2>`�3ڙ�����%��}��ϸ95�of���\��>=m�<�;tie��GB�uZv����a�]w���!=���Ϊ_>���K�ZMq-���#���5�u�˙���@�S=RI����V��%֨..���v<(�UK�Z�ݼ��uD+�q�A�ZcB��L2�Q���=;���}�Mq��=�ʠ2�H�m^�ފN1v4��w��<9��5����#) goaϧA��]�I���.�n�Ipd����1\ı\�:�Ŝ�@@��F����)ͬ^I�-����-%���aFO�s����i�5mK�i�?��\� �fhR��\��b\]�K��-KN�M�J03�x���~#��q��D�r��:���{�V/t�?H�K�9�Y�IAݑ���+M��[j�/�k���V�H��IE�Hۏ��-^�S��;�Y#�Q�HO��jn�q,�mf��,���j� ����+�Y���P��;q�P�M�׍�(�j&�q�\��;�%�?�&��b͓�ii,:kZG�[w��p{c��70��������Kk\O�Q������w� `�mR�Z��Y�e�}G��~+-��(�Y�T�Ez�+Q�+�񑏻QQ���ݻ����ݩ���9�d��O���B�v߉�U�kW)m�#�ڼ�]֭���uP�r :� ��+(�{�Ok7c��io�T��|�<����f�M^����RG���<�ǽ�./�-3�3���*�m���r���.�j�W�M��⩗f嘟��U%� �zb�M``�|��!ێ�ZD��ղ�)ߝ_�$b$�l;�A�;q���V0���p��ƈ� �$�0U�>��B�8u��^fJ��d�t����y���.���� �$���uWf9l�2h�}��E�SA�����k%��V�Z�Io)$�v�0��>�� *�d�;�ͨ&l�@$�+���g����{ymt���T~Y�径����0��e�6�ia����� c2y{	̐�9f_N{��:��y��i�l;��$��W��OPpOn�b���Nҥ}>YY.�h~����z�h������uw�%�Iy��3��}�>�k'��U�`nu�,n�@�P��`C8^ }��s�UQn׺�A���޼��dāA�{�`�?J���G:��i�j�Ы�pa=G�''4�Go�lt�k�ew{l��W8bCnc�u;f��P�;����܋ˤ2��J�8�3�$���I���\��g��]v�H��I�UTN{�c85�I��{�[���K�h���
����w�G�+���zm�B��9&+�rm��c��ޔSV	4�X����zv��J������>P���1����گ��V[�Vi�I
�L�� l��kKY�㼟S�������(0��)��|����Rk:�����i�qLb���a]�bw�2}:Uh�'m��sö�V�{o4��G^d1��;��<q��T�u;��;͆Q{�U�(T�����[ۛ��H�t�o����E FH�Ǡ���s^ v��c�Ғ�lA�w ~�lP�v���)��Le���Uy�J~e�q�kj���+�� a��w`\$XU#�>��U4�5��%�B-� �Fo��p�5���s��V���W!�:޿Ҫ�bM%�:j�P�5aq�C�Z��CԨ����X�Ϩ���ky&��rH�@����b�j�v�m�W�-,*т�!6��b�|4�:�mm���7��q۩�k!ݷ��%���O1�Q̳o'y ���S��g'?��'�הika&��,���lRr<�1^��*�S���A�?Ȭ���~�<Z���ngV��j$ �jd�fw?���!��omh��"�H��=*\dT.�s�I�B�wF��s����� �� �+���Fs	R� O�{�W��҄�y%�#�]7]���'������@��ח���ۊ;�TV՝�����%�:�p	��?�\ޖ[�M<�+"/�b�rGb��I�������
�Yז� 9�_�-b*Ł�HH��2{u&���To	-]��%;5С�O-�)�Fgn<t8?���ް�D�}�`�>TS������Ը�}U��`��������Vm����I�;������]�-�ަ�w ��q$~d0�2�����|g?�t�{�z�=��diH=�}J��I�[; ��rp�׎q^���E��z��i�	��q���ʺ�N˹�v����W�|i�o�b�7_�E{�@G~�����׊��O���?1����y�~�9k{���;k�] F�(2q��]:x�LԒ	l�ť��D�x���c��f�u����s(��h�,"��t�xݱՑ�?Jɹ�����<�/}p��A����������?�D��p����E�Lރj6��%��ŕ��$`��㷵u�ԵmrYov���l<�ρ��w8&��CGԙ�����d���F;�9�?�t���K���I�����e��^˷����t��ʄ�oS/�v��\�K��`4p��>\�<��W���Zd�u��&r��X��'����u�=Y���W�F����&:z�ϰ��N]_^f������G��}��Mەhs[B���d��unac&3� ��ʹMj����(SȷF!!k����{Qmi�L��6��[s��������췚������wh�`c=kD�;��3�X��ΞJ���Y	鏠������+f������o��Lՠ��]�,1:!R�
�{��T�K=$ژB]������-����yR|yjx�MZ�&��t�4V�<0�A������i��aG����]��]Iml��Ve��e�1��-���~d�kz�Ũ\�`��ܾ��ӵzǇ��3��3��K�'%�a\�_"�+4ڄĜ,��T^-��������#˅O;�rk�f�:`�Uٙ�H�0Gf� �F?ƸY$i��f'$�֖YY݋;�{�V`8^�Ҷ�TQ�Rm��=*�V�/<��	#�K����e������x{O�����((b%~Lq�z��MJ�;�f���2!��b��Q�n
y��h�Z�����H7yE����u�c�j��\����;X$,s���P9�݀�x�3[^�"-e+.'B·����=��T��+mJ���,ҙ�);����?�z
�mc�tsj6��X�� �s܁[�IuXUP�n�B�=��#ׯ��PZ��,�yo�*.�~q�-���8��js�bHI\�����A�
�QX,4ϲ�H�I2��r;/�����[O���F��o�B������Tw�a����L�30��f��Мs�5jWw�&����ό�y�<��MO}�{O�y��/�8�Ҡ�z�i�!N���ƣJ��x�W�����;��;�J{��<�&)�%�(y'��'�z����;���;��=��5��q��E�_oR�\���Ƶ���g��7��Gz�^؆��$�����������h-�rIȠ+��=Nr
��mb�X�`�����lD���8�=sX����R��c����X#6�ڢgq �v�L������Zɗ#��_��/�V��ɌI�y���F���E ӵM^��R��H��!-�ñR�8]���_O§�Αwơ��i���̱<��ݤ��n��ךy��/ͥۤI�[w�#݄��q�<S�k��ji���Ge)�!�q�1P\��I<;T�>�N���l�5�W�l�����ߎEii���<7���ILV�n r���<``�� Z�K�^�o!�%�_��I7�@�>�w�;�]Md��е7���!��~�q.��ˍ�#d����jӋ�vyc�F��m����u�����żǎv	�Ĳ�h��Xz��1\�������JSP�����bF w�=ɟcn��L��O��G��5�hh��á?^�ڳ�J�j1jy���@c�e����zu�Z�����]��̌|넑O�&2x������.� �'��ek��ڡq�w{c �}�it���6;�J�k�4U�&_�Obqǯ�i�|i���P��̐�6>��z��W�����)�JY`���\[C�2OR*
���CZ7��=f��(��(���8�u��S�V]{��/�H�1��A��Z��<>eK���_f�gv~x��U����ʱ, �T� �.�����1��.��W�ߜ�ϯj�����kWy�H�R7&z�޺_]�?
M� !G|?��<9���v����#rN����A�E���Ǐ.#���S��kޑ���v8�(���M���U��5eX0�ڳ�:��IY���rnn@ힵh��,��8�3����޴m-
���$ ��j'$�f��[���s�*#��<d� ��=+j�F>kL�Ԝ� X�U�ek=���i�����]�	���2 V{���ků�I���vIX��^%�%���U8Q�=��*��{��]�)f;ُˑ��շ4RO
�S�@�q�׷�[6����bH��p��Ð3�~��+r-7	B�?��1����L�\f�Տ��q޽���-�H�aQB��UM�N���0 QԌ}O��'�BOS�^�������QSY�"����v(��=�����}BMWV���;�$g9����+�׊�?��_,�=�Ӻ�׹�+�1�����j������58N3M@ �CO�M��m�����C��'�`\P��1<����?m��6&���v�Υ�������#��� "+���ki��G�ɀ�=k�Jҹn*I|�kwS���5��!�q�sYV�NETGo�kdԶ=;�k��{+-�;)gPx��Զv���!�mDh��3mQ��נ�����rnOB�����lN�
�d��lԚn�w{���,�~��q�sZ:Ɓ�����.��Wq������޲���ѧ�m�k�	ݺ/�� �
�$�"Qqvd���C����ds2¬>RF}� ư��In$i�$����+w@���U��D@���6��}:V<�F�z����lw �O��8��eJW�IZƴ�:���@�����V����uH��lf3�1�r��kwwV��k]��l�3ؕ�;g�z��mI!�#��p#A�=�De�vM��Bc�l>~���χ���p�"8^8&��
�Wօ�ՠ�� ��ի��4�}6�$q�q�� c�̬m
j�s�w�L�DJ@yF2N0+���E��}ٍN�޿�w� 5�0M�7->�� �ys�t��*���I��.�7��8��#Y���~�gi<����H�ں�l K�"� ,�8�@ϡ�*�+ls-uctK(�6��Č�r��3א{?:��6r�4��h��af���@ϩ${T���G�+���'�u�E8��k_\Y��Tǵ����� � ���a'�V0�"[y"�u��;4�&{��N*����'�n��n���w�q�a�8�G'=@����72�O2������H�*���u"�p!KO+ˎ63�㞽*U��zw:�/<~dQ1fWPD�2s����T���+V��D��.a��~�8�08�~�-muk��<������vc�8�;�V^�*H/����ڪs&��s� b�+[
�)�G�o��@�Pb��g
����ӿ֘%��(�<�C�y�,D����c�� ������2ʈ�6ڱ�O\�{���:�b�X��2H�D*�m�؃��Z�Y��Y�E�.�z��20Nr[� c�R�4���/�Z����� �)w*�y\o��� ����o>��x�� �+M]��=kN��(���}i�.����k��������'��z2����#�H3��
Xf��1��F����E8IIY�NwGU���F�y��k�i����H�_a�~��OJ�|)<w����XԢ���B����Oj�~������W�}��A�?]Eз�g<.���ǉ�O�:���M&��V,����<?t�]�dQ��6[���~�ͥ���mpډ+ �L��	=z�j��aK�
���_0���0rit�=#ӧ�m�;"R��������'���Sm,ʽ�љ�&�,t�b�P��L�G�($)�=�OÞ��"յ�n����FV\��#��~br@���{�P>&�o-#��)q$p�m�'��g�^:�����u��͕�ۤ�p�|����##��P����{����}[P��Ѭ�Ih�*»L�y2x��ӳ������9���y�%�{FT����<9k{,�WzS��F]�v�
x)�H5�o���]�j����ѦW�-ҀZ\u�9�u�U�ĥr�S���Lח�>b�l�s��%y���r����F���x����$T���8�?�nXGw���.���F�w:����u��t뎵��i�[\�a%��� �Z�sӐ;�翭J�B���cu>�me��"�>@S&g$c��O��W���x6�U�C��'�����v�NgKKk(lm���8e#�2�z�<�3ֳ����/o5'�i�as����=q�'��~·s�J�� ���I|���0=I�<b�|!�}���a���w��Ю5����P�?�u���k���X4�M���ǫ�zS��F���O����h�4�N��j���W��N�W4�.�$��k�#�jv� E��õr�t�eve^�3��F(�Fy�0
r6�M�N\��3��h�=1<�GC���XX�x�oC����B�4s/9�]>���c�B���� 
�M�tvS��i������6w���k&�Щ �3��x��#Y�/ �=�OE/���k��*3��O#5��G[�Ε'я�ҭ�9H�N1�f�"�P�v5TL�ǖuP�9c�V}����m�����?p�����S�('�Ir}Yе�P�]�(I8�_x���H���K��U�����r=+���\������f`���t w���k�է������:�e��{��eʟ+z�#�n�+K������3My���F,į$��&��ǘ>��j[{1sᛖ��f��r�Go֩�r�+��3.DjXя`:�mY>�XI��?̈�Ѯ�.88�A������bh.mt�l��S����J}���AY.�"����h�۫4�
�����c����%�t�2��O|p1�R���в��g ��j��#���� 99{���C���U��{gVb7+�ҳ[��3&L@�D�ڮ�8� ?Ұa�x'P����q0?&�Ns�Wao0��0��ҥ�Ӭux�]²/bG5JN�*
)�5{K��x����E)�y��
���� �V�),� �7����۶���^��M�kq	m8*J�*�7#�{�\��c����ټ2��w�>��=�Ji��b*Ǚ�^���-c�Ky=�RN軕�x}?ҶR�m+�Pٽ�rI)ށ9'wL���.����xv�L��ydg.Ҫ����m��Z�����q(�a���9��%gsf�M>&��v�u��pR4V��z�|�&�}S˙�a�y� W-����ז;{)P.�1��rs�=���<9�ã����7(��3i_CX�+�SJ+h����rzVN���w�-������9��&�]��dg�|/���O�!� ~����\���w�^6<�J�?,a��<�����>�{�^/�3�B<�����Es�L�I��b_;P���\������A �r7�kX�s�wv7tX�PY�^�<�X/.}�� 
�I�h0��ͮ�v'=�9�P�7O3B�C�3�=1����A�Z����s��$2������\�+�R�#��m������ڪ�w�8��*̚\�B�Oq@��'}���� c��@*�v6:bG<��	*[�F���ێO�=�7��$�K�o8����xS�Rx�}(���o��DIn���ʀ�u©�0s�j̒��oD#ϐ�(W$��������3�޼�x��H�ؑm��=Os�� +&��ɚ&Ti�]�L`��rO=1���p��{Zk�#��R/�bG9���$ѳf7R�K��,Qy��㏭Mz'��Y�dK����%~o��;s��WL�
=���F�F������یГ�qc-����~�&R���z����w?k��6�R�S�H3����Qק-an=�X����rF�,2EL6�Ğ6�����V����7�Ɨ��)�Eiu
���O)Dl�pU��x9��\��g� ���f�Cx��I"4����:��U|��v��?�Z�DF��Y�I�H�(�1Ɏ0C�pkW�� �j�I�0ew�[�����m���X�W�u�?1��%��y��J
�;:� ���[�S�P��m>�%C��WO��g�hL���1�)��,���q��J׺����Ź���_4L:��\�[w�?�j�N�ʚ��k�[���Y[NqdC1<7'�08���-��4�u�ޫG��a�\#�8�j������r[��kP9:f�"�{�Jg����ۨ21�����i��!�I�v���kkj���o�<mkhwM;�ޙ8�lb���<�Π����i���#kЏJ��u�}���l��G%�� ��9�8 �Z���S[M��P{�.I|���C�?O����D^�H%��sZ=�ܺ�2�e;Y_JʰG&œ���Wa�h�sG�l����@�c@�`�CךĴ���[�}&���K�G�+�I;�y g����֕ƻo��������~d�0�#��c�:�=lBM\��\A�j6:}���6 Iyg��ߌ1cМ��VLw���Ʈ�zZ�ɝf�}�L!ylz��J�d�Z��--���(.$��|�y'��>���\iڥ���߫Z�������\���z��u%�����>W(v���T�:;j�����ȏϝ+��ObҶ��gd����>��]X[m2�<�`�/П��)9��K�&���.�i���,�� �|e��a��XW�wS��k�%��<�K,��;ޙ�k�l�A�B7wb�R��E8�;�
�䰔S�M#�;�#�:?�1�ݱLqO\�ppGqI����/BX���̀I�K�\-��猎���'�#D��`GQZ�sϗ<��F���&Ϙ��Ь�C�ܑ�/sYN]�cdM���}�ڜ��q��]��}���Z���{��x���Å����Q��#�ԠѠc�6$a�G۟�ܼ֮il�BRH�q��Os\ؚ�6�����?=�$��S��Yt��$�� ��LSnt�>�^#+�˟1�p8�����%x�"E�3�L
u���ϐ!�(c#8ϯ� }+?n���ְv��4��Ռ�Ol����SˑO�듟ƬhZa���I�8 ���ۥ\���lƧf��2=Ϲ�s�RN�\C5�,�+��z�>���7�՝���]��v+�Cn��F��d<q�{�p1M�����#�O�@{� �z�'�ml�*���d��Oz���n��&<�&	+�t�O����ت���I6��,y�f2�̡V,)��;�k{�
܆���;`�OC�ά��QF��$*�Y��G��j�Q�i  )g ��S�tR���X�xzr�U���YkV��#p�V���ナ��{���Ll�6�Ât���3����~cַ�G�{h�Q�bz 2{�V^nP-�,�9!�k���e���J#��9�Z܋_�Q�unH� �v�u���$Kׁ������I�m��e��-FEm���{S���l���O�0ؿ�?�RM�rKvz<��$"�x���Y�"�K��%���
w�=��?1^s���X�բ��ɷ=b��{����9<�5j�s9T[D���wz��]_L��'s�z�V߅HK;�ß�s���ӿQ]G�@x/��ʙ�� �4ER���n������ ���c+�ǆUa�z�:z�t
g��Z������f��]�@-�}hm�;��;m0L&����r�Q����<rl�n�9�V)����� (�<�q�IAR���o9�T��͕�#}|�p3K��my�ߔ�Y���#;��9�y��k��_`7�[[Eg3'��g��t���!@�\��k1-�J�1H�Y�g'�P ��Ԍ¶<V��I�F�;��ۖ�3�n=��ֳn5id�ⲷ�Aʈ�A9Q��1�o���T����w{�����@d���U��@�Q����QX���{���-eU H#���e�h���6$�n��|"�z!9m�}���z
����!��cR1�
eʅ�ЁӞ)�����_�;K�6���?w���kw�Jd�H(������FyQ����)�g��lSk��Ǜ�A�=jψ#XmlQ|Ǻ`W
0���9��Z��V'����q������Ns��ߵ��܆x�� ��8�:1�Y�H,�d3L b�;� ��6��8Q���WU��u��j�m���o�=���]s�p~���O��Z�Ni+k"n{M��r�,�2���^G�)�1����1�������[E�g4�d�d��$-��NE^���-��Ws�A�OP?�u�~��n��l�év�Q��@F0������ǣ�HA�	(� ?���G��:і��eU�b��Z坜�u$�h6Ȅ���M&���>��6�^�����2���TJ�z2��=kG��<5���G4�����_�ҥ𮡣j�%�Ѱc!d%�`oS�B�C]$4�����R���U�-���0��\&�\3�]�ǆ"I�v�N�,�/���KC��m�夆dR��P�%�4^��m�پ�ko��c���<a�A��<�k:Uǈ�Ay�O+6� D
 � 
���䇍�U$#q���O}�CDk;���b~��t�W;{��ءk�{[_�n�3)�Zi��$�(�c�j/
��x�U�Y�F|�� �z�E{cco�L��G�;����M[V�9�WV}.�綱o�C� ) �g��e��Ftg��-� ��_^��c��>h�J���rG?���Er�z|^��d��F���O�� SU���͹7��~�l]��B��?�����h���"������ ����M�L��*������ߎ�qX,�����8��HJ��p�()*AEI è�O8���:�V"F$����ֵnڙ('���b�l�y�1���j��f#>L��kB����>�m&#z��. �`s�ϝ�c_g�8B���O����ww:�Z}Ɇ��)S=H�?
���?�8۠����	�?���tO�e�QG%��!�pRzб��@��z�5O �Zff�Q}n������ �O�M�NP�F��CwZ��E�+V�}��uV�E��Wz��r�;g��°��������s�� Uh���𵭶98,@�y� ?Z�-n���b��s<��͵KH�D�.���l�<�L�;�H��͜��W.Ȣ|�A��v���ϛvB�(L��3��y��*Y3����� eF�/ O3#o�x�J�E�+[��dU�N���O�1횳p�K#d�K ௷ኩr�	�ʅ�|��'vs�����:��Ô��gX�vv�N3����y��[Wq�4!O�� ���g��Ug)iiQa݈@HT�����34d@F�ǖ�̀��/� ���^rR[S���ڙv���h�M�Jv��'9>�枳Yi7
�K�I�99��֛ac<i,�$q���� �YS�n�p^B�7��=��5ؠ�ھ��R��F3����.��}��y �j>@;w�uR+�,�ڮ�m.�_�Ud�3A�  ��ql�I�]Q����y1R���wskTT���.���2:C��0��'����o��K�ۏ,��zg���b�j�V��Y>k�/�rd��S�ɥz̠a�#�֪+��A�l%+�d�c�mn�})ܑ�ړ�Z�v>�m��z��-Y�[�� g�RrHp��㉈WNH��u~�$�I'��3Ѓ�Ӛȱ�%�������� �žW�Мu�_��\��:!4s:�^]��zHH�y���o�M���Ь2�>�����5��PE������s���b��zV�w��EfwB��M[�)�{{�@ҤnO���#=�|qS}�5Ο",qH��d�2�|c��qY�N�#�!,��d�d�s� �����`<�%����F��g$dgw��[[X�2=r�Ηv�C5�v��
� ��{c����q�p���<eؼ`u��=*ˣ�7C"y��n�
,�t9�C�ֱ��3[,�w"�K�ȊK�q�DtqBM�~�j77V���+[�IHd�Y���翰��Q3:�-��"�|0p=��� ���z��.��,D�,�\+Hp3� zp9��˨%���m��y��ےG`��w������pђ�4/,ۏ���z���P��O:|��`K);�rO}��jоh.o-RG6����eʨ�1�ǩ�~���I��v'�V�,�!���Ϡ��ުKV&�gL��,��6@��}*	����p,�VDuf}�im��?�W�Cr�v����["Ų0�pO��ER�@����1Q��U��WS<6ײ1�e�(�ns�Һ�X�&����8�Z��"��"�� Ǖ�y{��?κMU��6��-�d`Nr�?�p;�z���MGImD+Gr�F� \ st�Ұ��9���+K۹���sO�R8?Һ�$��k9����t��S�H���K*�X�O�:� �����kaZ�!��>�����-�b�s�7��EQ𺥴I#m�m.6L�n��W(팄�Sq1���۹F����F���2�����~�q��h��i��v�I����})5[as������+/º����ձ:��I率�WA.!�/>��n�+g�[H��i1�� Yc`}G���zk��];�E(����8�^�"���nQ�֯�#7� ^��p�; �O4k���%c��:�O��#pK�����]�VS[�]�	iG(9��[Z��v���Y�E��r����M�)A�h���V)����7�b��Q;�º�g����V..���y���K��_�-l��s���6�[<��ҟ+z���Xۼ��$��SZڴRe�c��i]�H�q�GƓ�Dx�"�gx�F�'����j�6�2u��(4��߶��<��`��� �=x[�x����	�7�n��7����1[��Ԛȴ��Ub�82/m�_j������E�I�[�*D�WU2�!}�����=Fh��C(�(yVЃ]��Kr,���GvP�P�� ���bd����AB�A7ʮ��e�9���!$��p)4;���e!Rϖ�Us�V��lno��	�V���e���=���ˏ�I�4��)r������M���jϩ�zM�w0�ޫ0����Y��4;m�G+ H}����^k�k,��qhf����p���]���S.��K��d��dӎ��2RVgy�m᷸����	�}~��k_�P��,c��-v�>��Za��P/픕��T����?*����is��D(��m#c�$cڪ.��.�{�|;a�M���S�$���~_�mK��
�����`����V���_�R|�cl���'�#�5`��a*��B\�}�q׶x�*�e)s>�C�Ҍi�-l�4��4E���Ԟ�0?�s�Msyp�X� :|��5vYa���f�Dn '��s�:��T��U��D�->e+� �py�:P�O��V�m;�M�-�h��<�QQ>E=_��ȫ6�wr��0F���O��UL��Ie*��rw�5�u��р��Uu�s�\u��9��=��Z�4ܖ���n�bi<�Ȉ�M���O��_M	��tUS��N?>�-��\(�j�V-��{�~�:��zir��<n-�|�J˨�A��j������f��V�]�P�/A[4�9)�P�V�މ�C��৖ W<�ӶvM�F?�F��u� Ѕe���U������i��)c���S���(n�d>+��\g�^+N��W�`�s��E/�,`���jX�2n�����ֶ��8��j�_|�8�$�c��WG�o�.B$�TQ������X2�#/���z�Ŷ�whVO�s��J��oFt�?ds�62E4���H��!���	� Y�N牅� ������]l7���Z&��C�W7�r�>1� �5<ȗI���-�����ט�D��9�0�$�u@N��3�[i�W@�@���<�5��?c�e�yS�� ֭���#
�m]�:ޝm�a����K����Ϸ�h��8`Ya��IH�#fXc���zW���˙�Yq�8�$��<��w��$��g�$��G �B��'��V�[�ٝ��Ř��A��/(��`b/{�Ol��E������p,~Z�z��u<�]-����"�]Gs0��c;3�@������u,��Y>-��w��)#~��,0>�J��=BDOp��� b�l� ��#' �@���q)��Ih�"��Ep�B�� �'��z�./�..d���Y瀔�06��d�E��sU澸�K��q�bd�3�׎��Z���&݆[<�VBIe���\&D�_��� ~U��[�L$+G33���㏠�����;P�,�т����!G|�9�z��K7�(!���e-���s���u�5[\W����k��cV-��*;� ��&�j��K7 �[z�ݝ���$E�;|�V�r9�3Y�ro���%[��1��P´OM�z��2�2�/\���iO�俕�@���L���*�{F�e���[*�S̈́�0G�U�[�Okv�q,f;������
}��kFR$��JW�1��ֳnb��s��O�s���¸SG���\�6��,���ǐ�;��J��\ZɵD���E��6�� D��6�d=6��~�S<�r��
�.�0���2�"�E�)��-�
$�m���?�����k�иQax�f���?�WMB;˓�[��=����S��6�ȉ!��6q���U$���߅�|?�2�3Y�`�'�����m�خFNy�U~c����K�����_rwqԞ~���j�m����>��7X�kh�FG�އ�a�Hw��nNi]�
�J�R�-˙&bX���a}go��Yv�(<��zV-%�v�R�s���V����-���L�_kcr�N����S'.�?�n��ȫ�qҽ&-%tM*�9���T�0?�_Z��ĺt2�kP�"�@��x������3����8C��q��#�ʄ�H���ه��Ik?�eh�S�U8�ַ��Z%ޡ-�]�G��yݏҹ(�)�t�!f�`}Mk[�R�kv�Ip�҂ZE�('��Z-���wKB��nX��*��� �]U��w����G�5����s.��J��t��+�!������[�i��w�$������=�$�)�Nk��"�T���z���z��X�};+8;UGQ�Xm�d����_�h�jQ��L>l1�jz$B�w�s:�we�Mki��Q�S�aЊ�ĚN�����w�F��Y�u����9|�9P�r1�Ӑz��� j����B�bĆ������Z�s7Aѣ��i�e��G%��ջ�-F�G���b������r��ڻ�$)�rz��Ƒ.�~�Y��	#�L�tY��!�`���<
�h�Z�soҴ��ck�?�ƽ�m��bvƙl�+���q
��~��\i��py����$l�i�e��Ch�[ܢy�n���ޕ��\Zʱߔ�BrG�=��v�bx�L��~� ʸ����R�n�%�[W ;)��q���
�Ajz9~1�*2�M	�ˉ��,��k����}>��}*�������u$1�>��w`��B�E�xp1��ZMq�i����#+�z���?�՝H>k��Ur�����ӹ�Xm��;^���YĢ���&s���u��ѓs�	�Qߟn1�����s)]��c�����]72�j���d��&ٷ�y��4O)��d��>X���#9���H�J���Z����Z��,e���:�Gd�ش>M��)���G���'}�T�r�b���E�@��2�?�y?�O³�2rzR�#M3;uc�F~6��g=�wb���&󊎖� �lrd��AQ�ϽGo*r9��� �8�jMlzXL;܅co?s1��j]�G&;Xː98���H�۔;d(���Ix�;qx�vPt�����NJ笨ʕ94�q�m����2Lk�� �~���<v�K�������1ۘ�t��^F3�T�c�4�&t�lw4����t�MA)=�����(��0.�Ne���� �L�쭵+4��u1�7)�7p}+�ff{�~�|�tǭX�uc.�(}�t�+��s��DW-�0��S����5�#�:����O��jiw��дs�B��rKc��pqZw�Pj}����}��`yL���YN0x��ԑ�դ���:7S�6w�ȧʺ�$�� 8l��BGO^*x�m�l%�N�.�U ����׿5�ks�x��m+2�Q���s�֝�����2mR��R�~&��\Z�n4��nd��e1�DqE�l'�����򬉤6wr�d�&V04i�e��'�<���i�x}.]�_�����<��ps�4��B�� ȶ��B�{���Sӽ�kE���E�ۅ��:�a�}+�tD�����rޘ������ÄyZv�fX�PX�}�I�3Y���g�;E������@�0��^y���w���b��+t�J���S��=��ŭ���DXK�Y�mN:�:��?Y�'�����TtS��4C�jR3�?1���Z�ؒ;�+u' .x����d�`���w
]��x/�N��h��Y��H)I�u#���Q��.f	�P����������t��F��G����8�	)8�'��"�}�B�G����h�`RVܪ��O=~�����[�0��{lwc��C�����j�R-|��}M/����qP"�>�H�~tXz�@��/V�v� S����Vf�r�>py4���L�ro&i�*ŭ�ީ��8���nˍ�ǡ��1���;!7��<wx�������8=+?����t�������+ K��x�ۜ�޳��u�M�.�=<F2�������a������g�Rf�L}�NH8�kD��>�7�c����a�	�$�-��[�.���ɳ�+R�' mۂ�1\.���4��a�)�Y6Ww��K{;/�"Ğg`N?J��D7�=Ő[���f��EA���������&�]6.h��G$��|�s�{�G�����SL�31��}{V�n���%��7�����Y?b?Zk���6�m�������.܀ ��<����4mKMW�o& V5��!l��u����kr�$� ,8�+/l��`�BW�S�RI��2i;��|P4�C0i���p $� S^}q�mJ���ܴ�����Q���_i���n-�.�b�0U��rqϮ 5��4yR��� 㨢���m����TR	��s]L:Ŏ�cq���-e�G��`	���G��9.���H�`�g�r9�I�Zkɖ�_��l����D%v嗢�xSLT����S<������g�E�=M��$��߯�+GF��R��fb�3�����Q�Ɇ�X��$�����p�Kk#|ѯ�����V�$j%��ۡ�6�֘�D��ȸ��.�ɶ�~�����x�#�G���k���.��G�s����3�+�������wP�����?)l`���s�;�)7�_��;4���=ޏ�]B�$�)�����=H�ϥd�X5���!������N���P��Eĥ��� � t�V�����G;��tc�[������94��[����Β��4Q��}}=jy�e��
��6�yL�Q��ܰRa`s��������7kpҫ,���?&�����z��ޏg�z�)�`�w����s��ޱ���]�	9۞kF��m�$���B�Q�{��ɨle��B�m(f1��H�~�PR�^�V�F�H��� ��P��@o��ޖ�N�K&�!��[$�ҵ���6�GB����Aҳ�Mr��8&P�v1�G����=k8*���5���M�ݵk#:��df{�	zg����V��ݸT!N@�Gw}-䅤8�pV�Ĭx2�ՖÇBi*X�tgj,s@�i&�,Q�� ����xv�-�ߥL���
NsH�m#�=ȭmðM�`g��1��'��U�W	9�Th#ּ��n����(E&>8A���A�'�� ��.�[Ka �x�z}MOs8��2�)
�0=O�sYw�=̻�D�|����:q�w�]z��\V�kC�b�Ŝ���ԥ!�@Ub[��z��퍪 i�:��8�;�C[0iBf8Q�c��+Ug���(E]_��L���% L���Ko<��=�=�CmqvU�.䃹��,�l��F��O��u�i��
5#��'~�GT:\�[�c�=w{T���,�䔎W9#�Ec\��!I"�2�MV��q"�|��sZB��KC��V��97}�n���Б��ý(�P��9�����|�U��3�vh��~ky��`�?�g/u٘{7ʝ�dGs*I@ 8'#�z��e���V�!�)bK�pO��u��\�?J]�|ŗ<`��2kSJ,�uo��1o�����ݱ�>���N�HԵ�%x�3,x�����9�}� J�dl�z����	�a���)�V�����a�����!J�'E�{U������� >n-���V��Ɂ�c�3�~>Ec��i���5��!�(���V<�� �u	2�� `sQ���~b�W��Dz��9?�O�}�0�L_	�b�fr��6��mp�����R�'�*�q��O�YH�l�\�a�N���'��qMDQ��B{Ґ����5��D�A�~����aP^B�3��1#:(�v�=*�i�<99��0?:��H܁۞�О��׵���2hN*O<W�]�1���
��a��u�?�ZYV%bs��k������cjX����V�V��m�:;�V�W��Њh�����8�}��Y���<Me�NH�,X��d�����Rx:����#k��7��c��$���U/(q� �H=��������ɩD���S�L�q����-v���![$X�A*�?�^�滭H�4�)&���x�3>[z� &���o�J �y v�.�%es�o<Ye}�{9�[���@���k�����(�
;�|����5��=���oᨵ�����-���j8���j�P�$�	b(m�3���{=
�ҹ,��M^��V7m�YWv1�o��b�i�woi/��(���l�[�����"�3e��YI�y����םf�'�#����,�?J�Ki#�|5�D�0y,�e/�/RI=}N@�=�.���Igs|���x?Đi>�J2e�m����\�����Vڑ�������U7�ԫ7^Յ���\���Ġ������h^�R��YE���=:�s�i��:��0�(�S�	���V���?&��P�Y��9��?�u�VZ�#)��M|��ݟMAjW1�3t��?�x����z�����x�I鰁�s]Q���隄�}�i>�'@KF��Or:�\Ʒl�|z�)"��VI���H#�9�+�%�
rM+��)�F?x�֦��[����B��}��v\���-�f����;7j�&�"F�.��y,9��|6�p.5g[H�Ǖ��}GE?^}��M3@ҡ��[�y�q?�a);�tF�֧�� ��ܗA�l��K����zzW�=ƛ.!��pFR,VN��B��6^�
	���eUB��$�I�J��NjzWuu��x����pG� \zVUƏd��I��zU{d�oisx���_��r�mh��_U��*�ȉn�3�
�4�SWAgl��X�E$�@^�������j�]�����K�i����>R3Ҳu-&uS���1a@����@00>�V�	nw~��il<�5�僎:��� ʳ�?3���4��QZ���1+g@�=�.�<�����Tg���݄%�F�v���?�jι&�f%�`s�9g��J�R�]�:X�M%d�Cn�N�$n�c�.��>�GQ���A,̠�_w�*`��(E�$�=�U�f^������uӃN�`�V�+qz�cD_�m!*>�!�A��e����%�.���I4��r��#�KopVdX��O� ]j��{�n�JN��d:���(?z�g���OޤM>�$u� ����$:j$�����ZƟkxc|�In�����Uy�	Ej��;�D����(�ԞX�%VRy'ױ��ۏ�g��n���8>wr��`� �j���n��}�n���R���BB��<T�4���\c��XM^�A�);�#���"���3,L0�࿁�Ue�&HL��2c8S�����KI?� ����|t���ص��m�FNȬ`�jB��↥o���B;H�(�e���#:�Fhk�߳MX�_G����"<u*�pA+�S�֌�I�٭�n"T'<dsU���7˒=�1YbP;~����8�T���i�E�u~����_i� nOʡf=3&�P�c)Tw����?��Tт=��T^b�ƥBs���y�N��`��L��w'��T-ݱ�0(9<�Ri1�pTj�?L+~<Ud�G\� *�H�aq��;~��V��*��})�p9'��IC�1�9	���R�^� Η�N��n��%�2���}�3��V.Pd�%�]3S�ZYZ�$pK�1^���� 멀B9Zh�揞��4ǒ(�x���R�7� ��/��i�:��)�q�.>���ץK��Lw4����6�	��VF�I���V</��"��f�(��9�j�O�bG�K2F�&���:�}Kᶓq���'��E�I/txl�"B�W��҅+t%������<m鶚�:K��t?+u<�z�\߉�ϪdO-����5�C����^9�tm����~� ���qp�˷�c��hrW��A�f�v���D��V�I����u��5W�Ǉ4�ZK�AC�X,hG<��+�����G�ķK=*M;�k����SȂT��y���?"�<����ì�T&y8�A���Vz��M�Y(y���Q�|-�Kֺ{�6��J���S�g��xX�y<�4�v��Ƨ������e�'�;_�-Ŏc+�׍�=�?Z�\��f��y���� ����	o@?�ֱ<[��Od�s��܍!\)���Z��f�ʑ�9� ?Zʚ��e�9��f���b���w-	��B�@��{g�Q��S�V7�J\_J�yeV<�:
��+9���Z�g+�XDc,�ݡ��h��G�]����!v���5 c��irƜ����FJ����m�_�c����%~I<*�`+��������%�=ˏ�� �?_Sڲ<3}k�=��ą�};�����z~5�y�2���#��� ����&���])Ž	���H�h`#�x�O�R���KX�'�j�G&�!T�ь�� �����䍣$!B�x�^�kl�(�K�O�y�(+�qV�!T�ykrs�W7qq,�S�,@��xo���?�\U��l,���o��C'�����֥3�����.Ewg��0O�Ǩ��R�4k�@�H��B9�+����K�b9v��뜽�K���8X���s�r��C�þ�[�Q��b|�s�?1��"Kf���O�[��4q�I#:Ͽ�B��� �WE)���9I=
��Oc��a��?��"��KO�R�K�r��5�hd �m5��\N�x�Ԙ�U�z�ƶ�ס�ѝ��d��<��I����$�`V�0��y
V4���O%��![�QB�y�,V�;�z��>�����W!!VXS���� �:~B�'Q�>Ȝuw6��E��GK�,q�ȋ~Y>�� *ž�,����fG�?�u&��w"AbO�GB}}��g�J�Ws�z�J�QJR�z�f�(����g-pLsg��iB��$dU��E�8��U�����^��t�9��W���o��+����ƥ�R�	#�9#?�=�9nKO�[v���wf�"���9��KS�<�N0]��Ԓkh��Kp��<)�?�j��c��b�������N#,QT��&�	��Q��1��8]-wi)O��++���F�.�C��6����=j֭y��ۮp?O«�I�.�P͞�i��j��d�6����*���t�t���4{q�G$wǽR�1������Z��7�K����(l����������|�{��w,�%������NO�W/�(\��T�U�t�R���z����ְ�7$�pO5�����76��>��9���|��*����M{I�dt��~F!� �5jN.��QRVg�O���R� �U��:d7����|��� �W%wi-��9W��k��E4y�i8=6!�s��֓�J3Z\���]K8v�ON������-��=2�� Z��JX�D�7nH���LQl���@z�uc�'ܟ��m�[[�AS��R��R�{+W n�p��ǥ	�v�r���0b�Ķ﷞�� �*=��v}�����gU�K�������� ��$Ct�[�����~"�k��PH�ULC̍���jhqWG�����c���ǃM�����՝$,<��{K�G � 7Z҇�L���22�x��r�v���i��[�S��7C��U�闣[�c��?֡��)#���:\���W8Vw�:Њ�%,���� W�M��2�;hޟ��'��?��M&mkF���Bװ�(;yOaB�ch������O�g�'���Z�H�Q�ee�C��=�D�%�4	
3�YUF�T��6��Kȣϙ*�=H�&�d8��'޸9<]�� 1�� 5�ź���<�Z%'��=u;7'0��.*�O�
���^k���?ޞ�q�j�ͦ^�Eb8h���S�K2[]SGVg�do����Eד�f�n,�j˧j\��ʁ��}���I/���-&�3D�@���Tݧih=�u=}�4�B������j�=д���U��ꐟ1�O��{��F�Q��ˉÞ�HX~�*h��=�+�I�ߐ����jٔ�r��k?��&�`I�%�<����S_ռGr>�q,䟖%Q�Q�+Y�[���\��G���?i�5�"i�˱<��O�+T�wVR-Z�V����k[_6M���<�8�� ����c*C{pځ��f�m��L���q��\ӭU,%{��MAU�[���c��B'�;U���l��\����9��?<�Wm�!�tC�:Cokl�����~����s]&��;�_��Mo/�D��{�5��xf�C��b���w�����f����HE��.畗��
$�%�S��8�s=Nv�uWl��lr=�b�/�N�����BB�Y���`G��8�+n�a�� �[ׁ�۽c�h�M���6H���vƬw�'~�A���I&�y%��2�]�~_烎:���L�b8����ӎ�9��DR��X��#gv	�Os��Bܫ��hH�
A,FO�9�O=�*Ö� �r4x�g���#��)�V�y�c�t�6�p3��G������nY��,v�$�ݙv=y���X�ԧ�|��VB�lO�'#8�@���T���u$��1�s�g�ǽC}$F�ͅ����$�ק|~\b�<���Q(�C�@���u�h�jKR.����Y�A ������xm˴L��#J�=�g��Hն�#��@'$v?ε5]2$3��pO�%h.g��(F.M�yv��Au��ĶfFF�����OBG�tzn���Эŭ�W�(x��C��8${�u�}��l�p����T^F���*��O��Y�9j��ʪ;]�o�/� ��Y�$����{��R^�W�bH���e\�	�q��i��Ķw��lR��m��^�jί,Z�ϑ	���I!�� ���.K{o�ڞ"1���g�,C�$L��0O@?Ƨ�(a0���z��j�.�VX�.7�0���\���'�cH��W��jvr��}U,Tn��ɺQ$�D��Y��x�I��Uuzִ�m̂e�����N�1of�z�MtBkD�Z�ܯ6����@㖑� ��=��,�ƪ��=Ȫ��7����u�=�s4q2����'"�J�")K�NON�}���i%Y�T�>�E����9q؟AO�pۈc��j��l`kh+#��T枊����� UPr)lՊ� �ޜu���D�ĝ� T���I�a�RޖF��SRjȹnVXd���J���mz$��|����*��6���:b	:*�� "�C��Z^C7�/�v���ұN7ש�RnPӧW�;-5�xR�%��3�X/�nkd�q��8��V��ᱵ��F�0٫	"�A�o$�lr�n[�W2��Ea��=���d{�j�<��<���r�p߅K�2#!8�=1֩�[Ew�U���Z�{`�YcW��z�ք�d�&��GP�$�|��2xa�j�+��pQ�ea��֫gY�5�k�5���]�Y�D��ݾ`��"��m�$�� Н�=���U�W6�r�Hӵ[��T��q�e���� 
�ߩ���"��#�Kc��� =�SD&H� �1��t�����:�J��c9�R�oT���C��i	$:w<T����)I������>�:���� �m�����|O-�� ,7�a'�7�ǑX�j���� gl�f)��}j-f]B;��+ĒDGP:�ƚM=�����h�����6B����c����}5K�Y�/�#%O���O����s���eFW�����u�� �a�c���jR�a�����ԭta8J���%�嵍�����q��7���k��|K4��	gj��_(?_S\����w������K��1y��|�B� tV����̧%�}����d��[�ǥg5����v\�C�];E�p��.B��Ry��� HH�27�T }��y�**�)��VoC:���v8Aeq,�JHX`��ն�m�x. WUs�����9mgg��w���G~��i.#�,��ZG
�@�� �}���x�m:�`�7}�H�DLfB�6�>�?��?:ЏM���GR�|�`:�=~��d�o�I�S��d�{��ۊ-�nmw�cd����C��seBX�M����d��P�I�=�?_Z�,|K�j>M���&�\�R����,ء�휆� ��8Ϩ�j�h� �6�"ym\+�_�<g��ZR��;KU�ƶZ+>����x���I%?6���W����_�cg�&F����zע�wŲ�����q+�2�'P �Z~-����t�{�2��n��OC]~��zoNݏ.�9ҟ-O�<�Z��������� �=�1ڴ%�x�9 ������ʤf]�����sRkR-�-���4
�q�~��L�-fKڡe�V���$���J|���~�p��Cu�ȟk.x� �Zz�V��}���K(S?�r>������F�([{��$z����m�T"��w0 g8\����'�=�4S����]Ŧ麕�+Iq i�N8ϹL��BYg��,r	=k��զ�Ҭ,#Jq� �G�;S%�,��+�e#����ӊn�߸�t�]74t��mg)iW�}��}1߮MjCY� �F�f��1��8>����+:���Uq��;�g�;t��`�ee2�b�'������4�tb������	<��B�}�:7�f����_68K�F����� �}MZ��ڬn�qȱ#H�ݵNq��8�5RK;����Č��g����B��:4�"��a����?�A�
�,n<���`�����5�z��0k�L�<q�z��UBHZ��"Ć���r�oQ��Nj��W�ĺ�3#��q�   g��&�A(���CI'�� �z}rq�f�۱#��E$|����� :d��ʊ0��K(Q��~~��h���v�{=O��^�X�����A�V�u�� �J�I �ny'�+@so��4���i�9���U�ۏ�I���r#,HU�s\��۠T���e�+;c�a����<�ݎ��� ��Dbk��ڸ9��q��`�^!�[h>�̒`�������P����n�D��Ɨxd�:���O'��S�A�S{bt�*'��$�v_�:�� ��=�Ž�����u�
q�?SXQm�k�+��)�n-�k7̿C��һ[-F���r��#���m��L�'u�N=+wG�݌�HY'��,�G���r�Q�S����GC5��P��V#��\���_A#3G�o8Q-�����w3��w�$���q���޶���2wX�pg�QQ��R�7^���mu�y`��}�f��[�I��x�^��'R=�3Ueӭ&u2Z�e3��Nҹ2��7M����coo��2��j�֛w� �9\t�9�v��/ZGv��O�\���5�-�*���8�M�M�Ĩ�+�w(X`iX��U(���z��z]֑g��xܞ���qxkK�-U�~��~T��7�e6��Ko1��dK#���L�<��U����=<�#�UW����F�sSd���z��@� �J��n�eT�	�˨���w`j�����=� <�������5Xu��ɵ��}=j�G\��Q
g*?�v����6X�	^�qUK����cW<� �C/b*e�,P�ʎC���S1��M&z�B*���Ζ�l闖v%���Ȕi�LV�j2��X"��rEsWv�kKKFw/�� �8��I]F��@h� ��Z7��+�aՔ:)B�n>���󔻽��b�� ����ŵ�<�qؚ�[�mn��y�/&�$e� �%+;��i>F���8�[�ţ[	6�!�Ԟ?�ݫOY��5+K�H�Ii�`2}��*�υm�飶fE�n���E��!��F1��B�Q�N�Z)���I+�4�;��
mE�L��H�d�?��==O5���Bi��<����V��\��I{ 	!�p#A��
�%��nrOS�h��z�j�m�u{ &[��r�ǀ+�Ӽ2!��pB�'�NZ����7Ăq�3ӟ�� �WQm�&1#!�Q�zW'�$6;0�E�=Y��V�v]���=�kB�<@��de' �[���5Ţ��,1e��~�b���68����^_5�g�eml��f�d�W���76����Qc��-&:`�'��{՛�c;B��~p22�Β��m+̄HUI������}�D�̛崱�e��A1���� � �z�N�wM����J<�`�� �	���a�6jڳ��9��+t�1������lZ�2�2�*��l��ps]�tӽ̔ڛV/I:[�ᦝ���QTm�{RKt��vǻr��S�9�:w��2mF� %�ú4����� ��U5B#{h�ώWU�26���u'���Dav�rI;8t���eX]]]Q[$����ޣ�u��+iWP[�nx.��X��o�ð8<~>��]�X�y�"V1p����?"s��k�<���U�`I`1��a�}��+Zu'NJHέ(U�����W��� �4��ь�����?�y.�o$�m��x����r�{υu3}m&�xC�a�é�2==��~"xh�wĲ"-g>dG��^�9ei.��V��zr�~C46-N;��|,1m �Nz~�|#7��S�h�@�;�y�@ ~5�=̰ۘHѻ�㎟�ih�B���]���T�*��n��r� �:����l�ZZ�Vs�vK�=�e��}�i����N=�l�ܫ�£lj�����γwDU��:S791��;���=���McS]��)e
>nwp{��d[HЇyTJb"@�y��~2j����И����:�g�r?,{Vv2.��A����p�`��tOP�G}2�eܤ���nq���L�ͷ� D~���@$����x��i�̻X�ѫ��R8����up���k�%>�����z�9���6g�@�N��d��@ z�犋S�͟���E����p����Es��?�D��"9;$������VЅ�lM�$��a�Į�r�=:~��yp�����w1�U�?G�Wue��̈�N��}�#�q�̕�nc-���vT�1ִ��}��ע+g����C� ��>��s�j�E�a#����� �$w��/ڛ�U|�h���:�s�b�j��VaC��$汜9�k
*��<sP�Bv�X��,��	��5��#M��%�'$�sV<Ew���M����>Á������t�k
J��Z�I����v�#ҷ�.�u{�I�q���j���_����q��O:� g_�q�G��6��M,ҹ�G�A�y��a��g��G���w�4�ɆQ�&�i@�d*ޑ(�M������V�A��ւ�ˑG�ț��nk��ۡЕ����mk�C���<�vȫ�{����iɩ�N��w.A<�޹�7F�������U�F�=>����Ma��% ��� ��ПC�R��i=��q-���ڻ��ge������G�e�V���s(88��N�����X�Il��Ƀ¿N}2*/�֒���7�����!��S����g5��-�>.>�>�r;�p��P_��aYi���_�'���	=�� �J϶���M���f[�#��8 v�*�d�4u�ϯ�q�B��rA^����T��D���>}����v�>��O� 	�-ݢG�o�M.VW�GF�9�y�A.9�� J�_[��<r�$|����lv����.B��POf����}��.�9�8�{�|�������(���m=j��'��؊�tU�,>�� �U�����5�&2s��Ry�xrG�^�b7�T��c4�4g�ʷL��� ��G5�� ���hM�!�'�u�L���껆F%X��3�>�E�t��sg��r\L�&�^K^@̏�z��� :�G�n-'�o��:�ޕ�6�&�-�����Vѕ��۩i��Db˞�,O��V\`��,*��ʓ�\�r`~��_��Ȫ6��	��P��Z�n!���Ж
;�� 
���ҭ�`$I|E�� ���_ƶ��&��~Ixbz=Ƹ_j"�X���a�Fe
qL�fс��na�qZ^����9`71��ҹ���=Nk�|3m���KA ���St�+n���U����6�
�r0�iU���R4�&P�dʨS�����zƆG��'� ��J$X��QA�Rv����ws��ۈ���f`���Z��1����0A1 0y�����RH�#��I�����0?q�7�����6�q��N*�WЎ8���`9S����g"�q"���-Ia�w�#=��V���B�FI^�����_ΰ�$�)W�o��}�O����q��`��ٙrm�Uui!'�x�I�x��QOs�.Q�����A��q��v��B{���F�&�8UN�^rGoa֥�x�Q�,�����2Os�ֻ�;Z����TiI�[�d��nwی�?�z��yy,���I�K�Y����..oZIOͷq�>��U�,�7�$�1����N�ؙվ�ċ2	Qr@�Ĝ�A�AֵFك��&_ ���V<a����#RK"�����=z�Zq�+�Z5H�B*��#��s��Jʤt4��k���O�m�w�0#O(xَ����C�E]S��H�0�5��!�`˗`ð88�+���߁��w�Z%q�8�?#]X)�.�<�Ɲ���g�A��*�S<`�N��a6�2��z7*�A^��G��&�@�9<�c�^b�C($�r�+ �#Ҧ��s�����D�twgS����̭������>�+T\�6�s2��aJ?P;{9��\�WC�M��Ӏ_Jݷ�W6�+d�.����m�"��#˺<yl�r��׸#�J��D��%ʬRITC�.3�R{w�b"�U@<�A9|zzv�=�Pڴ�Cp��W�R��v�?���Ͽ~�����E-�U
0̤�����=z�U�q�yo�˱\�N�� J�Q����%@
F �@Gn��nO��!h��+9�8���U���sz'�m��G��A�Ą�]�y���֥���D���1����3�W�����m��<c#�w�m%�һ;��b���_ް�y�lWI��a��.s���ס����ޘ�V�I��p����quli��N�\������Qvv/r�1,ē�NI�qK<�(�!?(Q�j晡˨��&;e8yH� ���k�]��"��0�Y��?�V���naJ��3�,�����UF�(�$}�٦O���\1�c��R�� }���Ԯ/[2���G T	|��5��ճ��l��7�g9FP�vj��q�m�tGV�N����$�/��kOM����2��u+�g� �Q9R�����
r�^�/�K�s�zT�}u�q����V��Z�`�wܹ��d���P��Kyr_D�L~F^}��x��(�(�6�Ʈ�D�h�-VP2�3�f���)�h%�Q���?�I�xg�":�Ҧ@9 c?�t��m^4S'<��8J�^�R�N�lt���&�i{<H^�4\oS��:��WV���V��6o*�A� �$v��R6<��������Rq�����}j�f����"f����܍����� �Y�g[?N��[�?�|#Wf�}CI���~�u{��E��}�,��sn�d���}��vFj��9�J�Ĉ2�kc���j�ز:�xϙ?��Z�c��_���Ҳ#��)��9�5t�*u,�/M�FYc������j��}4Q��Y\�k��G�y��7��ǘ�w���l�-����?�S~����;O\.D�$�������5�i �<�L� *�d
�;T���� Wu��U��J�������� ӌ�F#�ڹ^�Xj�n瀏�p#�����U�����zw�/��eE����A�U�?��� }�*�JK�J�_SN��;}N��p���v\Ex���އ��W�~�� ]O����>��� �i�Y�q��>U���{v�d��<��_ޠ���G����1���bw���j�� "�%f;��!����f���x���W<c�5�R��rkCC� �^�� \�� B��� �+O�)$\vl϶]�(��,2kԴ��UX"��`=�ym��|�z�����ʹs)4�ו�/�7�B���O~��Z�:E��� ��}N}�l��� ��jb�ԟ���˶��уn6���X#d �<�Ϝ�.�
ؚ�6��݆;�ԒǕ��ƥ_�� ���R{0]\��2��2r:��k��l��J�Y�9���ӶkzO������aj_���_�
ָme�WH��@�I)*A�6~��늊젎@�#"��?���S����z�G��OO�����F/Nc��BgyJ@�,s/LB�{
�ŶUl��ď�TZ���"� �q� *�>��� Ыd�FW՗V,��;8�$�s���Y9%a�2fUR?�r8�+_���������� v���oE�cu�����������+��ݛ��f&)FA<�GC��z�!� �4��]�����?��j���a���gl,�a�B��b?�c
�$� �@����צ�G�Ո��st��D�rݬΙ�[
���Z��nLgF��@�?�r/�]d� y� �cTh��v�$�h���1�~��-�G=�++Jg�n
9!I��+f/�����\�� �ş�p?��Anl�i�
�Y��<��=�x���h���`��� ��i���}[�#��G}�  k���*�q4O6ebp	��Z�_xN+[h��	f�T�1����V���� ���W��������$��B)���mv�Y���S��?Os)#N�" ����}��=�z���_���kʹ���� �F�쎮T��c[T��DFމ���6�I$���Ӛ�j�HƤ�<=��F{⺽3C>lf���H[��Ƴ���v���]���n?�y��D����%���4�.�-��:n���=I��mg���QWq9�7���M?�A�����+C� ���­Zm��SԌ"��)ǾU}�mRsǷ��:�^�ZK[u�	��Xu�ܞ����5��� ��o�觇��5�ME�?�RQu
əF̟�p�t��z����y�k�t��U5�q�  �?��<U� #}������t������Сs���gj�2y\�`��GR����� �a����W��X� ���#]�zҨڑ�Zj���ǒ�<�� �W-G��L����vȠ�� �V��|AV$� U'�[7���*�.��-ј�	�����[�۝��Z����Y7��'ֺi�˩����j���FG٪�3Z���2��Q��zWG�o�s�W5�� �^�����T�<�fOrJ!�.T��³�M�T�	�*�}�� �-Te����LP�d�(oOJ|_y~��U��A�~T�ք���WUi� P�5�T(��